`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:54:05 12/14/2016 
// Design Name: 
// Module Name:    MC14495_ZJU 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MC14495_ZJU(D0, 
                   D1, 
                   D2, 
                   D3, 
                   LE, 
                   point, 
                   a, 
                   b, 
                   c, 
                   d, 
                   e, 
                   f, 
                   g, 
                   p);

    input D0;
    input D1;
    input D2;
    input D3;
    input LE;
    input point;
   output a;
   output b;
   output c;
   output d;
   output e;
   output f;
   output g;
   output p;
   
   wire XLXN_5;
   wire XLXN_10;
   wire XLXN_14;
   wire XLXN_19;
   wire XLXN_37;
   wire XLXN_38;
   wire XLXN_39;
   wire XLXN_40;
   wire XLXN_41;
   wire XLXN_42;
   wire XLXN_43;
   wire XLXN_45;
   wire XLXN_46;
   wire XLXN_47;
   wire XLXN_48;
   wire XLXN_49;
   wire XLXN_50;
   wire XLXN_51;
   wire XLXN_52;
   wire XLXN_55;
   wire XLXN_56;
   wire XLXN_57;
   wire XLXN_58;
   wire XLXN_59;
   wire XLXN_60;
   wire XLXN_61;
   wire XLXN_62;
   wire XLXN_63;
   wire XLXN_64;
   wire XLXN_65;
   wire XLXN_66;
   wire XLXN_67;
   
   AND4  XLXI_1 (.I0(XLXN_19), 
                .I1(XLXN_14), 
                .I2(D2), 
                .I3(D3), 
                .O(XLXN_60));
   AND4  XLXI_3 (.I0(D0), 
                .I1(D1), 
                .I2(D2), 
                .I3(XLXN_5), 
                .O(XLXN_59));
   AND3  XLXI_4 (.I0(XLXN_14), 
                .I1(XLXN_10), 
                .I2(XLXN_5), 
                .O(XLXN_58));
   AND3  XLXI_5 (.I0(D0), 
                .I1(D1), 
                .I2(XLXN_5), 
                .O(XLXN_57));
   AND3  XLXI_6 (.I0(D1), 
                .I1(XLXN_10), 
                .I2(XLXN_5), 
                .O(XLXN_56));
   AND3  XLXI_7 (.I0(D0), 
                .I1(XLXN_10), 
                .I2(XLXN_5), 
                .O(XLXN_55));
   AND3  XLXI_8 (.I0(D0), 
                .I1(XLXN_14), 
                .I2(XLXN_10), 
                .O(XLXN_52));
   AND3  XLXI_9 (.I0(XLXN_14), 
                .I1(D2), 
                .I2(XLXN_5), 
                .O(XLXN_51));
   AND2  XLXI_10 (.I0(D0), 
                 .I1(XLXN_5), 
                 .O(XLXN_50));
   AND4  XLXI_11 (.I0(XLXN_19), 
                 .I1(D1), 
                 .I2(XLXN_10), 
                 .I3(D3), 
                 .O(XLXN_49));
   AND3  XLXI_12 (.I0(D0), 
                 .I1(D1), 
                 .I2(D2), 
                 .O(XLXN_48));
   AND3  XLXI_13 (.I0(D1), 
                 .I1(D2), 
                 .I2(D3), 
                 .O(XLXN_45));
   AND4  XLXI_14 (.I0(XLXN_19), 
                 .I1(D1), 
                 .I2(XLXN_10), 
                 .I3(XLXN_5), 
                 .O(XLXN_43));
   AND3  XLXI_15 (.I0(D0), 
                 .I1(D1), 
                 .I2(D3), 
                 .O(XLXN_42));
   AND3  XLXI_16 (.I0(XLXN_19), 
                 .I1(D2), 
                 .I2(D3), 
                 .O(XLXN_41));
   AND3  XLXI_17 (.I0(XLXN_19), 
                 .I1(D1), 
                 .I2(D2), 
                 .O(XLXN_40));
   AND4  XLXI_18 (.I0(D0), 
                 .I1(XLXN_14), 
                 .I2(D2), 
                 .I3(XLXN_5), 
                 .O(XLXN_39));
   AND4  XLXI_19 (.I0(D0), 
                 .I1(D1), 
                 .I2(XLXN_10), 
                 .I3(D3), 
                 .O(XLXN_38));
   AND4  XLXI_20 (.I0(D0), 
                 .I1(XLXN_14), 
                 .I2(D2), 
                 .I3(D3), 
                 .O(XLXN_37));
   AND4  XLXI_21 (.I0(XLXN_19), 
                 .I1(XLXN_14), 
                 .I2(D2), 
                 .I3(XLXN_5), 
                 .O(XLXN_47));
   AND4  XLXI_22 (.I0(D0), 
                 .I1(XLXN_10), 
                 .I2(XLXN_14), 
                 .I3(XLXN_5), 
                 .O(XLXN_46));
   INV  XLXI_23 (.I(D3), 
                .O(XLXN_5));
   INV  XLXI_26 (.I(D2), 
                .O(XLXN_10));
   INV  XLXI_27 (.I(D1), 
                .O(XLXN_14));
   INV  XLXI_28 (.I(D0), 
                .O(XLXN_19));
   OR4  XLXI_29 (.I0(XLXN_38), 
                .I1(XLXN_37), 
                .I2(XLXN_47), 
                .I3(XLXN_46), 
                .O(XLXN_61));
   OR4  XLXI_30 (.I0(XLXN_42), 
                .I1(XLXN_41), 
                .I2(XLXN_40), 
                .I3(XLXN_39), 
                .O(XLXN_62));
   OR3  XLXI_31 (.I0(XLXN_45), 
                .I1(XLXN_43), 
                .I2(XLXN_41), 
                .O(XLXN_63));
   OR4  XLXI_33 (.I0(XLXN_49), 
                .I1(XLXN_48), 
                .I2(XLXN_47), 
                .I3(XLXN_46), 
                .O(XLXN_64));
   OR3  XLXI_34 (.I0(XLXN_52), 
                .I1(XLXN_51), 
                .I2(XLXN_50), 
                .O(XLXN_65));
   OR4  XLXI_35 (.I0(XLXN_57), 
                .I1(XLXN_56), 
                .I2(XLXN_55), 
                .I3(XLXN_37), 
                .O(XLXN_66));
   OR3  XLXI_36 (.I0(XLXN_60), 
                .I1(XLXN_59), 
                .I2(XLXN_58), 
                .O(XLXN_67));
   OR2  XLXI_37 (.I0(LE), 
                .I1(XLXN_61), 
                .O(a));
   OR2  XLXI_38 (.I0(LE), 
                .I1(XLXN_62), 
                .O(b));
   OR2  XLXI_39 (.I0(LE), 
                .I1(XLXN_63), 
                .O(c));
   OR2  XLXI_40 (.I0(LE), 
                .I1(XLXN_64), 
                .O(d));
   OR2  XLXI_41 (.I0(LE), 
                .I1(XLXN_65), 
                .O(e));
   OR2  XLXI_42 (.I0(LE), 
                .I1(XLXN_66), 
                .O(f));
   OR2  XLXI_43 (.I0(LE), 
                .I1(XLXN_67), 
                .O(g));
   INV  XLXI_44 (.I(point), 
                .O(p));
endmodule

